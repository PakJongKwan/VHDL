--COUNT_8BIT.VHD
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY COUNT_8BIT IS
PORT(
	RESETN : IN STD_LOGIC;   	--RESET
	CLK : IN STD_LOGIC;	--CLOCK BUTTON
	
	COUNT_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)	--LED OUTPUT
);
END COUNT_8BIT;
ARCHITECTURE HB OF COUNT_8BIT IS
SIGNAL CNT_8BIT : STD_LOGIC_VECTOR(7 DOWNTO 0);
BEGIN
PROCESS(RESETN, CLK)
BEGIN
	IF	RESETN = '0' THEN
		CNT_8BIT <= (OTHERS => '0');
	ELSIF CLK'EVENT AND CLK='1' THEN
		IF CNT_8BIT="11111111" THEN 
			CNT_8BIT <= (OTHERS => '0');
		ELSE
			CNT_8BIT <= CNT_8BIT + 1;
		END IF; 
	END IF;
END PROCESS;
COUNT_OUT <= CNT_8BIT;
END HB;
